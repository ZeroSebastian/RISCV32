	component riscv_system is
		port (
			clk_clk           : in  std_logic                     := 'X';             -- clk
			const_high_export : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			leds_export       : out std_logic_vector(7 downto 0);                     -- export
			reset_reset_n     : in  std_logic                     := 'X';             -- reset_n
			switches_export   : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component riscv_system;

	u0 : component riscv_system
		port map (
			clk_clk           => CONNECTED_TO_clk_clk,           --        clk.clk
			const_high_export => CONNECTED_TO_const_high_export, -- const_high.export
			leds_export       => CONNECTED_TO_leds_export,       --       leds.export
			reset_reset_n     => CONNECTED_TO_reset_reset_n,     --      reset.reset_n
			switches_export   => CONNECTED_TO_switches_export    --   switches.export
		);

